----------------------------------//1.dataflow modeling//---------------------------------------------
module half_adder(
                 input a,b,
		 output sum,carry
		);
   assign sum=a ^ b;
   assign carry=a & b;
endmodule

---------------------------//2.gate-level_modeling//---------------------------------------------------
module half_adder(input a,b,
                  output sum,carry);
  
  xor w1(sum,a,b);
  and x1(carry,a,b);
endmodule
------------------------------------//3.behavioural modeling//----------------------------------------
module half_adder(input a, b,
                  output reg sum,carry);
  
  always@(*) begin
    sum=a^b;
    carry=a&b;
  end
endmodule

----------------------------------------------------//4.modeling using the switchcase//
module half_adder(input a,b,
                  output reg sum,carry);
  always@(*) begin
    case({a,b})
      2'b00:
      begin
        sum=0;carry=0;
      end
      2'b01:
      begin
        sum=1;carry=0;
      end
      2'b10:
        begin
          sum=1;carry=0;
        end
      2'b11:
        begin
          sum=0;carry=1;
        end
    endcase
  end
endmodule 
----------------------------------------------//5.functional level_modeling//--------------------------------------------------------------------------
module half_adder(input a,b,
                  output sum,carry);
  
  function[1:0]half_adder;
    input a,b;
    begin
      half_adder[0]=a^b;
      half_adder[1]=a&b;
    end
  endfunction
  assign {carry,sum}=half_adder(a,b);
endmodule

-----------------------------------------//6.structural modeling//-------------------------------------------------------------------------------
module half_adder(input a,b,
                  output sum,carry);  
wire don1,don2,don3;
  
  not t1(not_a,a);
  not t2(not_b,b);
  and a1(don1,not_a,b);
  and a2(don2,a,not_b);
  xor x1(sum,don1,don2);
  and e1(carry,a,b);
endmodule
   
-------------------------------------//7.parameter_initialization _method//--------------------------------------------------------------------------
module half_adder#(
  		parameter Width=1
)(input[Width-1:0] a,b,
  output [Width-1:0]sum,carry);
  
  assign sum=a^b;
  assign carry=a&b;
endmodule

--------------------------------------//8.look_up_table_method//----------------------------------------------------------------------------------------
module half_adder(input a,b,
                  output reg sum,carry);
  always@(*)begin
    case({a,b})
      2'b00:{sum,carry}=2'b00;
      2'b01:{sum,carry}=2'b10;
      2'b10:{sum,carry}=2'b10;
      2'b11:{sum,carry}=2'b01;
    endcase
  end
endmodule

---------------------------------------//9.using generated block//----------------------------------------------------------------------


module halfadder(input a,b,
                 output sum,carry);
 genvar i;
 generate 
   for (i=0;i<1;i=i+1)begin:sub_half
      assign sum=a^b;
      assign carry=a&b;
    end
  endgenerate
endmodule
  
